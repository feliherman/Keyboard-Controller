library ieee;
use ieee.std_logic_1164.all;

entity Decoder is
	port(Cod:in std_logic;
	Intrare:in std_logic_vector(0 to 7);
	Iesire:out std_logic_vector(0 to 6));
end entity;

architecture A_Decoder of Decoder is 	 
signal A,B:std_logic_vector(0 to 6);
begin 

	with Intrare select
	
	A <= "0000010" when "00011100",   --a
	"1100000" when "00110010",		    --b
	"1110010" when "00100001",		    --c
	"1000010" when "00100011",			--d
	"0010000" when "00100100", 		--e
	"0111000" when "00101011",			--f   
	"0000100" when "00110100",			--g
	"1101000" when "00110011",			--h
	"1001111" when "01000011",			--i
	"0000011" when "00111011",			--j
	"1111000" when "01000010",			--k
	"1111001" when "01001011",			--l
	"0110000" when "00111010",			--m
	"1101010" when "00110001",			--n
	"1100010" when "01000100",			--o
	"0011000" when "01001101",		   --p
	"0010100" when "00010101",			--q
	"1111010" when "00101101",      	--r	
	"0100100" when "00011011",			--s
	"1001110" when "00101100",			--t  
	"1100011" when "00111100",			--u
	"1011100" when "00101010",			--v
	"0000110" when "00011101",			--w
	"0110110" when "00100010",			--x
	"1000100" when "00110101",			--y
	"0010010" when "00011010",			--z
	"0000001" when "01000101",			--0
	"1001111" when "00010110",			--1
	"0010010" when "00011110",			--2
	"0000110" when "00100110",			--3
	"1001100" when "00100101",			--4
	"0100100" when "00101110",			--5
	"0100000" when "00110110",			--6
	"0001111" when "00111101",			--7
	"0000000" when "00111110",			--8
	"0000100" when "01000110",		 	--9
	
	"1110111" when "01011000",       -- CapsLock

	"0111111" when "11100000",     --E0  <--,-->
	"0111111" when "01101011",     --6B
	"0111111" when "01110100",     --74
	"0111111" when "11110000",     --F0

	"1111111" when others;	
	
	
	     with Intrare select
	
	B <= "0001000" when "00011100",     --A
	"0000000" when "00110010",				--B
	"0110001" when "00100001",          --C
	"0000001" when "00100011",          --D	
	"0110000" when "00100100",          --E
	"0111000" when "00101011",          --F
	"0100001" when "00110100",          --G
	"1001000" when "00110011",          --H
	"1001111" when "01000011",          --I
	"1000011" when "00111011",          --J
	"0110100" when "01000010",          --K
	"1110001" when "01001011",          --L
	"0010101" when "00111010",          --M
	"0001001" when "00110001",          --N
	"0000001" when "01000100",          --O
	"0011000" when "01001101",          --P
	"0010100" when "00010101",          --Q
	"0010000" when "00101101",			   --R
	"0100100" when "00011011",          --S
	"0001111" when "00101100",          --T
	"1000001" when "00111100",          --U
	"1010101" when "00101010",          --V
	"0100011" when "00011101",          --W
	"1001000" when "00100010",          --X
	"1001100" when "00110101",          --Y
	"0010010" when "00011010",          --Z 
	"0000001" when "01000101",				--0
	"1001111" when "00010110",				--1
	"0010010" when "00011110",				--2
	"0000110" when "00100110",				--3
	"1001100" when "00100101",				--4
	"0100100" when "00101110",				--5
	"0100000" when "00110110",				--6
	"0001111" when "00111101",				--7
	"0000000" when "00111110",				--8
	"0000100" when "01000110",			 	--9
	
	"1110111" when "01011000",    	   -- CapsLock
	
	  --PT CODURILE SAGETILOR AVEM NISTE VALORI OARECARE
	"0111111" when "11100000",  	   --E0  <--,-->
	"0111111" when "01101011",  		--6B
	"0111111" when "01110100",     	--74
	"0111111" when "11110000",     	--F0
		
	
	"1111111" when others;
	
	
	  with Cod select		--DACA E SCRIS MARE SAU MIC
	 Iesire <=B when '1',
    A when others;	
	
end architecture;